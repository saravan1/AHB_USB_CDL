// $Id: $
// File name:   ahb_lite_usb.sv
// Created:     4/21/2021
// Author:      Lohith Chittineni
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: AHB USB Top Level Design

module ahb_lite_usb
(
    input wire clk,
    input wire n_rst,
    input wire dplus_in,
    input wire dminus_in,
    input wire haddr,
    input wire hsel,
    input wire 

);



endmodule
